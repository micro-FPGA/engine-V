module ROM512K16 (clk,	addr, dout);
input clk;
input [8:0] addr;
output [15:0] dout;
reg [15:0] dout; 
reg [8:0] addr_r; 

always @(posedge clk)  begin : process_clk  addr_r <= addr; end

always @(addr_r) begin : process case (addr_r)

  0 : begin dout <= 16'h E0D0; end
  1 : begin dout <= 16'h 2E0D; end
  2 : begin dout <= 16'h EFDF; end
  3 : begin dout <= 16'h 2E1D; end
  4 : begin dout <= 16'h 2D70; end
  5 : begin dout <= 16'h B818; end
  6 : begin dout <= 16'h BA00; end
  7 : begin dout <= 16'h B808; end
  8 : begin dout <= 16'h EA4B; end
  9 : begin dout <= 16'h E0D0; end
  10 : begin dout <= 16'h BB48; end
  11 : begin dout <= 16'h BA10; end
  12 : begin dout <= 16'h 0F44; end
  13 : begin dout <= 16'h BA00; end
  14 : begin dout <= 16'h 19D1; end
  15 : begin dout <= 16'h FFD3; end
  16 : begin dout <= 16'h CFF9; end
  17 : begin dout <= 16'h B818; end
  18 : begin dout <= 16'h E043; end
  19 : begin dout <= 16'h E052; end
  20 : begin dout <= 16'h B808; end
  21 : begin dout <= 16'h EFEC; end
  22 : begin dout <= 16'h EFFF; end
  23 : begin dout <= 16'h E0D0; end
  24 : begin dout <= 16'h B368; end
  25 : begin dout <= 16'h 7061; end
  26 : begin dout <= 16'h 0F77; end
  27 : begin dout <= 16'h 2B76; end
  28 : begin dout <= 16'h BB48; end
  29 : begin dout <= 16'h BA10; end
  30 : begin dout <= 16'h 0F55; end
  31 : begin dout <= 16'h 1F44; end
  32 : begin dout <= 16'h BA00; end
  33 : begin dout <= 16'h 19D1; end
  34 : begin dout <= 16'h FFD3; end
  35 : begin dout <= 16'h CFF4; end
  36 : begin dout <= 16'h 8370; end
  37 : begin dout <= 16'h 5FEF; end
  38 : begin dout <= 16'h 09F1; end
  39 : begin dout <= 16'h FDF6; end
  40 : begin dout <= 16'h CFEE; end
  41 : begin dout <= 16'h FFF7; end
  42 : begin dout <= 16'h CFEC; end
  43 : begin dout <= 16'h B818; end
  44 : begin dout <= 16'h 2CA0; end
  45 : begin dout <= 16'h 2CB0; end
  46 : begin dout <= 16'h C027; end
  47 : begin dout <= 16'h E0D4; end
  48 : begin dout <= 16'h C001; end
  49 : begin dout <= 16'h E0D6; end
  50 : begin dout <= 16'h 2CCA; end
  51 : begin dout <= 16'h 2CDB; end
  52 : begin dout <= 16'h 2EAE; end
  53 : begin dout <= 16'h 2EBF; end
  54 : begin dout <= 16'h C014; end
  55 : begin dout <= 16'h E040; end
  56 : begin dout <= 16'h E050; end
  57 : begin dout <= 16'h E060; end
  58 : begin dout <= 16'h E070; end
  59 : begin dout <= 16'h 2FE1; end
  60 : begin dout <= 16'h 95E2; end
  61 : begin dout <= 16'h 7FE0; end
  62 : begin dout <= 16'h FD07; end
  63 : begin dout <= 16'h 60E8; end
  64 : begin dout <= 16'h 23EE; end
  65 : begin dout <= 16'h F029; end
  66 : begin dout <= 16'h EFF1; end
  67 : begin dout <= 16'h 8340; end
  68 : begin dout <= 16'h 8351; end
  69 : begin dout <= 16'h 8362; end
  70 : begin dout <= 16'h 8373; end
  71 : begin dout <= 16'h 2DDA; end
  72 : begin dout <= 16'h FFD1; end
  73 : begin dout <= 16'h C009; end
  74 : begin dout <= 16'h E0D0; end
  75 : begin dout <= 16'h EFF2; end
  76 : begin dout <= 16'h E3E0; end
  77 : begin dout <= 16'h 82A0; end
  78 : begin dout <= 16'h 82B1; end
  79 : begin dout <= 16'h E1E0; end
  80 : begin dout <= 16'h 82C0; end
  81 : begin dout <= 16'h 82D1; end
  82 : begin dout <= 16'h C0CF; end
  83 : begin dout <= 16'h E0D4; end
  84 : begin dout <= 16'h 0EAD; end
  85 : begin dout <= 16'h 1CB0; end
  86 : begin dout <= 16'h 2CCA; end
  87 : begin dout <= 16'h 2CDB; end
  88 : begin dout <= 16'h 2DEA; end
  89 : begin dout <= 16'h 2DFB; end
  90 : begin dout <= 16'h 8100; end
  91 : begin dout <= 16'h 8111; end
  92 : begin dout <= 16'h 8122; end
  93 : begin dout <= 16'h 8133; end
  94 : begin dout <= 16'h FD02; end
  95 : begin dout <= 16'h C172; end
  96 : begin dout <= 16'h 2FE2; end
  97 : begin dout <= 16'h 95E2; end
  98 : begin dout <= 16'h 7FE0; end
  99 : begin dout <= 16'h FD17; end
  100 : begin dout <= 16'h 60E8; end
  101 : begin dout <= 16'h EFF1; end
  102 : begin dout <= 16'h 80C0; end
  103 : begin dout <= 16'h 80D1; end
  104 : begin dout <= 16'h 80E2; end
  105 : begin dout <= 16'h 80F3; end
  106 : begin dout <= 16'h FD05; end
  107 : begin dout <= 16'h C097; end
  108 : begin dout <= 16'h EF7F; end
  109 : begin dout <= 16'h EF6F; end
  110 : begin dout <= 16'h 2F42; end
  111 : begin dout <= 16'h 9542; end
  112 : begin dout <= 16'h 704F; end
  113 : begin dout <= 16'h 9532; end
  114 : begin dout <= 16'h 2F53; end
  115 : begin dout <= 16'h 6F50; end
  116 : begin dout <= 16'h 7F30; end
  117 : begin dout <= 16'h 2B43; end
  118 : begin dout <= 16'h FD53; end
  119 : begin dout <= 16'h C003; end
  120 : begin dout <= 16'h 705F; end
  121 : begin dout <= 16'h E060; end
  122 : begin dout <= 16'h E070; end
  123 : begin dout <= 16'h FF04; end
  124 : begin dout <= 16'h C054; end
  125 : begin dout <= 16'h FD16; end
  126 : begin dout <= 16'h C009; end
  127 : begin dout <= 16'h FD15; end
  128 : begin dout <= 16'h C043; end
  129 : begin dout <= 16'h FD14; end
  130 : begin dout <= 16'h C01B; end
  131 : begin dout <= 16'h 0D4C; end
  132 : begin dout <= 16'h 1D5D; end
  133 : begin dout <= 16'h 1D6E; end
  134 : begin dout <= 16'h 1D7F; end
  135 : begin dout <= 16'h CFB3; end
  136 : begin dout <= 16'h FD15; end
  137 : begin dout <= 16'h C007; end
  138 : begin dout <= 16'h FD14; end
  139 : begin dout <= 16'h C026; end
  140 : begin dout <= 16'h 254C; end
  141 : begin dout <= 16'h 255D; end
  142 : begin dout <= 16'h 256E; end
  143 : begin dout <= 16'h 257F; end
  144 : begin dout <= 16'h CFAA; end
  145 : begin dout <= 16'h FD14; end
  146 : begin dout <= 16'h C005; end
  147 : begin dout <= 16'h 294C; end
  148 : begin dout <= 16'h 295D; end
  149 : begin dout <= 16'h 296E; end
  150 : begin dout <= 16'h 297F; end
  151 : begin dout <= 16'h CFA3; end
  152 : begin dout <= 16'h 214C; end
  153 : begin dout <= 16'h 215D; end
  154 : begin dout <= 16'h 216E; end
  155 : begin dout <= 16'h 217F; end
  156 : begin dout <= 16'h CF9E; end
  157 : begin dout <= 16'h 2F48; end
  158 : begin dout <= 16'h 714F; end
  159 : begin dout <= 16'h F031; end
  160 : begin dout <= 16'h 0CCC; end
  161 : begin dout <= 16'h 1CDD; end
  162 : begin dout <= 16'h 1CEE; end
  163 : begin dout <= 16'h 1CFF; end
  164 : begin dout <= 16'h 0D41; end
  165 : begin dout <= 16'h F7D1; end
  166 : begin dout <= 16'h 2D4C; end
  167 : begin dout <= 16'h 2D5D; end
  168 : begin dout <= 16'h 2D6E; end
  169 : begin dout <= 16'h 2D7F; end
  170 : begin dout <= 16'h CF90; end
  171 : begin dout <= 16'h FD15; end
  172 : begin dout <= 16'h CFE4; end
  173 : begin dout <= 16'h FF14; end
  174 : begin dout <= 16'h CFDD; end
  175 : begin dout <= 16'h 2F48; end
  176 : begin dout <= 16'h 2F53; end
  177 : begin dout <= 16'h 9552; end
  178 : begin dout <= 16'h 714F; end
  179 : begin dout <= 16'h F391; end
  180 : begin dout <= 16'h FF52; end
  181 : begin dout <= 16'h C007; end
  182 : begin dout <= 16'h 94F5; end
  183 : begin dout <= 16'h 94E7; end
  184 : begin dout <= 16'h 94D7; end
  185 : begin dout <= 16'h 94C7; end
  186 : begin dout <= 16'h 0D41; end
  187 : begin dout <= 16'h F7D1; end
  188 : begin dout <= 16'h CFE9; end
  189 : begin dout <= 16'h 94F6; end
  190 : begin dout <= 16'h 94E7; end
  191 : begin dout <= 16'h 94D7; end
  192 : begin dout <= 16'h 94C7; end
  193 : begin dout <= 16'h 0D41; end
  194 : begin dout <= 16'h F7D1; end
  195 : begin dout <= 16'h CFE2; end
  196 : begin dout <= 16'h FD14; end
  197 : begin dout <= 16'h C003; end
  198 : begin dout <= 16'h E8D0; end
  199 : begin dout <= 16'h 0EFD; end
  200 : begin dout <= 16'h 0F7D; end
  201 : begin dout <= 16'h 1AC4; end
  202 : begin dout <= 16'h 0AD5; end
  203 : begin dout <= 16'h 0AE6; end
  204 : begin dout <= 16'h 0AF7; end
  205 : begin dout <= 16'h F008; end
  206 : begin dout <= 16'h CF68; end
  207 : begin dout <= 16'h E041; end
  208 : begin dout <= 16'h CF67; end
  209 : begin dout <= 16'h FF06; end
  210 : begin dout <= 16'h C00F; end
  211 : begin dout <= 16'h 0EC4; end
  212 : begin dout <= 16'h 1ED5; end
  213 : begin dout <= 16'h E0D4; end
  214 : begin dout <= 16'h 0EAD; end
  215 : begin dout <= 16'h 1CB0; end
  216 : begin dout <= 16'h 2D4A; end
  217 : begin dout <= 16'h 2D5B; end
  218 : begin dout <= 16'h EFDE; end
  219 : begin dout <= 16'h 22CD; end
  220 : begin dout <= 16'h 2CAC; end
  221 : begin dout <= 16'h 2CBD; end
  222 : begin dout <= 16'h E0D4; end
  223 : begin dout <= 16'h 1AAD; end
  224 : begin dout <= 16'h 08B0; end
  225 : begin dout <= 16'h CF57; end
  226 : begin dout <= 16'h 2DEC; end
  227 : begin dout <= 16'h 2DFD; end
  228 : begin dout <= 16'h 0FE4; end
  229 : begin dout <= 16'h 1FF5; end
  230 : begin dout <= 16'h 8140; end
  231 : begin dout <= 16'h FD14; end
  232 : begin dout <= 16'h C014; end
  233 : begin dout <= 16'h FD15; end
  234 : begin dout <= 16'h C00A; end
  235 : begin dout <= 16'h FD16; end
  236 : begin dout <= 16'h CF4B; end
  237 : begin dout <= 16'h FF47; end
  238 : begin dout <= 16'h CF49; end
  239 : begin dout <= 16'h EF5F; end
  240 : begin dout <= 16'h FF57; end
  241 : begin dout <= 16'h CF47; end
  242 : begin dout <= 16'h EF6F; end
  243 : begin dout <= 16'h EF7F; end
  244 : begin dout <= 16'h CF46; end
  245 : begin dout <= 16'h FDE0; end
  246 : begin dout <= 16'h CF38; end
  247 : begin dout <= 16'h FDE1; end
  248 : begin dout <= 16'h CF36; end
  249 : begin dout <= 16'h 8151; end
  250 : begin dout <= 16'h 8162; end
  251 : begin dout <= 16'h 8173; end
  252 : begin dout <= 16'h CF3E; end
  253 : begin dout <= 16'h FDE0; end
  254 : begin dout <= 16'h CF30; end
  255 : begin dout <= 16'h 8151; end
  256 : begin dout <= 16'h FF16; end
  257 : begin dout <= 16'h CFEE; end
  258 : begin dout <= 16'h CF36; end
  259 : begin dout <= 16'h FF06; end
  260 : begin dout <= 16'h C04E; end
  261 : begin dout <= 16'h FD04; end
  262 : begin dout <= 16'h C005; end
  263 : begin dout <= 16'h FD03; end
  264 : begin dout <= 16'h C04A; end
  265 : begin dout <= 16'h FF02; end
  266 : begin dout <= 16'h C048; end
  267 : begin dout <= 16'h CF60; end
  268 : begin dout <= 16'h EFF2; end
  269 : begin dout <= 16'h E1E0; end
  270 : begin dout <= 16'h E0C0; end
  271 : begin dout <= 16'h 2FD1; end
  272 : begin dout <= 16'h 77D0; end
  273 : begin dout <= 16'h 23DD; end
  274 : begin dout <= 16'h F4A9; end
  275 : begin dout <= 16'h FF34; end
  276 : begin dout <= 16'h C003; end
  277 : begin dout <= 16'h FD35; end
  278 : begin dout <= 16'h C00E; end
  279 : begin dout <= 16'h E8C0; end
  280 : begin dout <= 16'h 82A0; end
  281 : begin dout <= 16'h 82B1; end
  282 : begin dout <= 16'h E0D3; end
  283 : begin dout <= 16'h FF24; end
  284 : begin dout <= 16'h 60D8; end
  285 : begin dout <= 16'h 23CC; end
  286 : begin dout <= 16'h F009; end
  287 : begin dout <= 16'h E0D7; end
  288 : begin dout <= 16'h E2E3; end
  289 : begin dout <= 16'h 83C0; end
  290 : begin dout <= 16'h E2E0; end
  291 : begin dout <= 16'h 83D0; end
  292 : begin dout <= 16'h E5E0; end
  293 : begin dout <= 16'h 80A0; end
  294 : begin dout <= 16'h 80B1; end
  295 : begin dout <= 16'h CF2E; end
  296 : begin dout <= 16'h 2FE2; end
  297 : begin dout <= 16'h 7FE0; end
  298 : begin dout <= 16'h FF37; end
  299 : begin dout <= 16'h C001; end
  300 : begin dout <= 16'h 60E4; end
  301 : begin dout <= 16'h 8140; end
  302 : begin dout <= 16'h 8151; end
  303 : begin dout <= 16'h 8162; end
  304 : begin dout <= 16'h 8173; end
  305 : begin dout <= 16'h FF16; end
  306 : begin dout <= 16'h C009; end
  307 : begin dout <= 16'h 2EC2; end
  308 : begin dout <= 16'h E0DF; end
  309 : begin dout <= 16'h 22CD; end
  310 : begin dout <= 16'h 0CCC; end
  311 : begin dout <= 16'h FD17; end
  312 : begin dout <= 16'h 18C1; end
  313 : begin dout <= 16'h 24DD; end
  314 : begin dout <= 16'h 24EE; end
  315 : begin dout <= 16'h 24FF; end
  316 : begin dout <= 16'h FF15; end
  317 : begin dout <= 16'h C010; end
  318 : begin dout <= 16'h FD14; end
  319 : begin dout <= 16'h C005; end
  320 : begin dout <= 16'h 2AC4; end
  321 : begin dout <= 16'h 2AD5; end
  322 : begin dout <= 16'h 2AE6; end
  323 : begin dout <= 16'h 2AF7; end
  324 : begin dout <= 16'h C009; end
  325 : begin dout <= 16'h EFDF; end
  326 : begin dout <= 16'h 26CD; end
  327 : begin dout <= 16'h 26DD; end
  328 : begin dout <= 16'h 26ED; end
  329 : begin dout <= 16'h 26FD; end
  330 : begin dout <= 16'h 22C4; end
  331 : begin dout <= 16'h 22D5; end
  332 : begin dout <= 16'h 22E6; end
  333 : begin dout <= 16'h 22F7; end
  334 : begin dout <= 16'h 82F3; end
  335 : begin dout <= 16'h 82E2; end
  336 : begin dout <= 16'h 82D1; end
  337 : begin dout <= 16'h 82C0; end
  338 : begin dout <= 16'h CEE8; end
  339 : begin dout <= 16'h FD06; end
  340 : begin dout <= 16'h C012; end
  341 : begin dout <= 16'h FD04; end
  342 : begin dout <= 16'h C010; end
  343 : begin dout <= 16'h 2F41; end
  344 : begin dout <= 16'h 0F44; end
  345 : begin dout <= 16'h 714E; end
  346 : begin dout <= 16'h FD07; end
  347 : begin dout <= 16'h 6041; end
  348 : begin dout <= 16'h 2FD3; end
  349 : begin dout <= 16'h 95D2; end
  350 : begin dout <= 16'h 7ED0; end
  351 : begin dout <= 16'h 2B4D; end
  352 : begin dout <= 16'h 2F53; end
  353 : begin dout <= 16'h 9552; end
  354 : begin dout <= 16'h 7057; end
  355 : begin dout <= 16'h FD37; end
  356 : begin dout <= 16'h 6F58; end
  357 : begin dout <= 16'h 0EC4; end
  358 : begin dout <= 16'h 1ED5; end
  359 : begin dout <= 16'h 2FE2; end
  360 : begin dout <= 16'h 95E6; end
  361 : begin dout <= 16'h FD30; end
  362 : begin dout <= 16'h 68E0; end
  363 : begin dout <= 16'h 7FE8; end
  364 : begin dout <= 16'h EFF1; end
  365 : begin dout <= 16'h 8180; end
  366 : begin dout <= 16'h 8191; end
  367 : begin dout <= 16'h 81A2; end
  368 : begin dout <= 16'h 81B3; end
  369 : begin dout <= 16'h FF06; end
  370 : begin dout <= 16'h C02A; end
  371 : begin dout <= 16'h FD15; end
  372 : begin dout <= 16'h C003; end
  373 : begin dout <= 16'h E8D0; end
  374 : begin dout <= 16'h 26FD; end
  375 : begin dout <= 16'h 27BD; end
  376 : begin dout <= 16'h 1AC8; end
  377 : begin dout <= 16'h 0AD9; end
  378 : begin dout <= 16'h 0AEA; end
  379 : begin dout <= 16'h 0AFB; end
  380 : begin dout <= 16'h FF16; end
  381 : begin dout <= 16'h C016; end
  382 : begin dout <= 16'h FD14; end
  383 : begin dout <= 16'h C002; end
  384 : begin dout <= 16'h F010; end
  385 : begin dout <= 16'h CEC5; end
  386 : begin dout <= 16'h F0B8; end
  387 : begin dout <= 16'h 0F11; end
  388 : begin dout <= 16'h 711E; end
  389 : begin dout <= 16'h 9532; end
  390 : begin dout <= 16'h 2FD3; end
  391 : begin dout <= 16'h 7ED0; end
  392 : begin dout <= 16'h 2B1D; end
  393 : begin dout <= 16'h 703F; end
  394 : begin dout <= 16'h FD33; end
  395 : begin dout <= 16'h 6130; end
  396 : begin dout <= 16'h 7137; end
  397 : begin dout <= 16'h FD07; end
  398 : begin dout <= 16'h 6038; end
  399 : begin dout <= 16'h FD34; end
  400 : begin dout <= 16'h 6E30; end
  401 : begin dout <= 16'h 0EA1; end
  402 : begin dout <= 16'h 1EB3; end
  403 : begin dout <= 16'h CEC2; end
  404 : begin dout <= 16'h 28CD; end
  405 : begin dout <= 16'h 28CE; end
  406 : begin dout <= 16'h 28CF; end
  407 : begin dout <= 16'h FF14; end
  408 : begin dout <= 16'h C002; end
  409 : begin dout <= 16'h F749; end
  410 : begin dout <= 16'h CEAC; end
  411 : begin dout <= 16'h F339; end
  412 : begin dout <= 16'h CEAA; end
  413 : begin dout <= 16'h FF04; end
  414 : begin dout <= 16'h C011; end
  415 : begin dout <= 16'h 2F48; end
  416 : begin dout <= 16'h 2F59; end
  417 : begin dout <= 16'h 2F6A; end
  418 : begin dout <= 16'h 2F7B; end
  419 : begin dout <= 16'h FD16; end
  420 : begin dout <= 16'h CF06; end
  421 : begin dout <= 16'h FD15; end
  422 : begin dout <= 16'h CF1D; end
  423 : begin dout <= 16'h FD14; end
  424 : begin dout <= 16'h CEF4; end
  425 : begin dout <= 16'h FF36; end
  426 : begin dout <= 16'h CED8; end
  427 : begin dout <= 16'h 1AC8; end
  428 : begin dout <= 16'h 0AD9; end
  429 : begin dout <= 16'h 0AEA; end
  430 : begin dout <= 16'h 0AFB; end
  431 : begin dout <= 16'h CEF6; end
  432 : begin dout <= 16'h 2DEC; end
  433 : begin dout <= 16'h 2DFD; end
  434 : begin dout <= 16'h FD14; end
  435 : begin dout <= 16'h C013; end
  436 : begin dout <= 16'h FD15; end
  437 : begin dout <= 16'h C011; end
  438 : begin dout <= 16'h 8380; end
  439 : begin dout <= 16'h FFF7; end
  440 : begin dout <= 16'h C00D; end
  441 : begin dout <= 16'h FDF5; end
  442 : begin dout <= 16'h C00B; end
  443 : begin dout <= 16'h E0CA; end
  444 : begin dout <= 16'h B800; end
  445 : begin dout <= 16'h E4DD; end
  446 : begin dout <= 16'h 0DD1; end
  447 : begin dout <= 16'h F7F1; end
  448 : begin dout <= 16'h B980; end
  449 : begin dout <= 16'h 9587; end
  450 : begin dout <= 16'h 6880; end
  451 : begin dout <= 16'h 0DC1; end
  452 : begin dout <= 16'h F7C1; end
  453 : begin dout <= 16'h CE81; end
  454 : begin dout <= 16'h CE80; end
  455 : begin dout <= 16'h FDE0; end
  456 : begin dout <= 16'h CE68; end
  457 : begin dout <= 16'h FD14; end
  458 : begin dout <= 16'h C004; end
  459 : begin dout <= 16'h FDE1; end
  460 : begin dout <= 16'h CE64; end
  461 : begin dout <= 16'h 83B3; end
  462 : begin dout <= 16'h 83A2; end
  463 : begin dout <= 16'h 8380; end
  464 : begin dout <= 16'h 8391; end
  465 : begin dout <= 16'h CE75; end
  466 : begin dout <= 16'h FD04; end
  467 : begin dout <= 16'h C01D; end
  468 : begin dout <= 16'h FF05; end
  469 : begin dout <= 16'h CE71; end
  470 : begin dout <= 16'h FF03; end
  471 : begin dout <= 16'h CE88; end
  472 : begin dout <= 16'h 9532; end
  473 : begin dout <= 16'h 7F37; end
  474 : begin dout <= 16'h FD24; end
  475 : begin dout <= 16'h 6038; end
  476 : begin dout <= 16'h 9522; end
  477 : begin dout <= 16'h 702E; end
  478 : begin dout <= 16'h 2EC3; end
  479 : begin dout <= 16'h EFD0; end
  480 : begin dout <= 16'h 22CD; end
  481 : begin dout <= 16'h 2AC2; end
  482 : begin dout <= 16'h 2ED1; end
  483 : begin dout <= 16'h 22DD; end
  484 : begin dout <= 16'h 703F; end
  485 : begin dout <= 16'h 2AD3; end
  486 : begin dout <= 16'h E0D4; end
  487 : begin dout <= 16'h 0EAD; end
  488 : begin dout <= 16'h 1CB0; end
  489 : begin dout <= 16'h 2D4A; end
  490 : begin dout <= 16'h 2D5B; end
  491 : begin dout <= 16'h 0CAC; end
  492 : begin dout <= 16'h 1CBD; end
  493 : begin dout <= 16'h E0D8; end
  494 : begin dout <= 16'h 1AAD; end
  495 : begin dout <= 16'h 08B0; end
  496 : begin dout <= 16'h CE48; end
  497 : begin dout <= 16'h 2F73; end
  498 : begin dout <= 16'h 2F62; end
  499 : begin dout <= 16'h 2F51; end
  500 : begin dout <= 16'h 7F50; end
  501 : begin dout <= 16'h E040; end
  502 : begin dout <= 16'h FD05; end
  503 : begin dout <= 16'h CE43; end
  504 : begin dout <= 16'h 2D4A; end
  505 : begin dout <= 16'h 0D5B; end
  506 : begin dout <= 16'h CE40; end
  507 : begin dout <= 16'h CE4B; end
 default: begin dout <= 16'h xxxx; end
endcase
end

endmodule
